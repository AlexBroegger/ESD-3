library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity txtest is
    port(
        clk :in std_logic

    );
end txtest;