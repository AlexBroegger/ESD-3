library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UART is
    port(
        clk :in std_logic


    );
end UART;

