library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rxtest is
    port(
        clk :in std_logic

    );
end rxtest;